library IEEE;
use IEEE.STD_LOGIC_1164.ALL;



entity Not32TB is
Port ( );
end Not32TB;

architecture Behavioral of Not32TB is

begin


end Behavioral;
